module and_t (input a, input b, output y);
  assign y = a & b;
endmodule